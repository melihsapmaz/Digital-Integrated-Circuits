* SPICE3 file created from inverter.ext - technology: scmos

.option scale=0.12u
.include ./tsmc025.lib

Vdd VDD 0 2.5
Vin A 0 PULSE(0, 2.5, 0ns, 10ns, 10ns, 20ns, 40ns)
CL Y 0 1fF
.TRAN 1ns 100ns

M1000 Y A GND Gnd nfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1001 Y A VDD Vdd pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
C0 Y A 0.04fF
C1 VDD Y 0.28fF
C2 GND Y 0.16fF
C3 GND Gnd 0.18fF
C4 Y Gnd 0.29fF
C5 A Gnd 0.69fF
C6 VDD Gnd 0.20fF