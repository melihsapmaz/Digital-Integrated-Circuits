magic
tech scmos
timestamp 1732306995
<< ntransistor >>
rect -5 -41 -3 -31
rect 3 -41 5 -31
rect 27 -41 29 -31
rect 35 -41 37 -31
rect 62 -41 64 -31
rect 70 -41 72 -31
rect 102 -41 104 -31
rect 110 -41 112 -31
rect 143 -41 145 -31
rect 151 -41 153 -31
rect 177 -41 179 -31
rect 185 -41 187 -31
rect 215 -41 217 -31
rect 223 -41 225 -31
rect 253 -41 255 -31
rect 261 -41 263 -31
rect 287 -41 289 -31
rect 295 -41 297 -31
rect 338 -41 340 -31
rect 346 -41 348 -31
rect 370 -41 372 -31
rect 378 -41 380 -31
rect 405 -41 407 -31
rect 413 -41 415 -31
rect 445 -41 447 -31
rect 453 -41 455 -31
rect 486 -41 488 -31
rect 494 -41 496 -31
rect 520 -41 522 -31
rect 528 -41 530 -31
rect 558 -41 560 -31
rect 566 -41 568 -31
rect 596 -41 598 -31
rect 604 -41 606 -31
rect 630 -41 632 -31
rect 638 -41 640 -31
<< ptransistor >>
rect -5 21 -3 41
rect 3 21 5 41
rect 27 21 29 41
rect 35 21 37 41
rect 62 21 64 41
rect 70 21 72 41
rect 102 21 104 41
rect 110 21 112 41
rect 143 21 145 41
rect 151 21 153 41
rect 177 21 179 41
rect 185 21 187 41
rect 215 21 217 41
rect 223 21 225 41
rect 253 21 255 41
rect 261 21 263 41
rect 287 21 289 41
rect 295 21 297 41
rect 338 21 340 41
rect 346 21 348 41
rect 370 21 372 41
rect 378 21 380 41
rect 405 21 407 41
rect 413 21 415 41
rect 445 21 447 41
rect 453 21 455 41
rect 486 21 488 41
rect 494 21 496 41
rect 520 21 522 41
rect 528 21 530 41
rect 558 21 560 41
rect 566 21 568 41
rect 596 21 598 41
rect 604 21 606 41
rect 630 21 632 41
rect 638 21 640 41
<< ndiffusion >>
rect -6 -41 -5 -31
rect -3 -41 3 -31
rect 5 -41 6 -31
rect 26 -41 27 -31
rect 29 -41 35 -31
rect 37 -41 38 -31
rect 61 -41 62 -31
rect 64 -41 70 -31
rect 72 -41 73 -31
rect 101 -41 102 -31
rect 104 -41 110 -31
rect 112 -41 113 -31
rect 142 -41 143 -31
rect 145 -41 151 -31
rect 153 -41 154 -31
rect 176 -41 177 -31
rect 179 -41 185 -31
rect 187 -41 188 -31
rect 214 -41 215 -31
rect 217 -41 223 -31
rect 225 -41 226 -31
rect 252 -41 253 -31
rect 255 -41 261 -31
rect 263 -41 264 -31
rect 286 -41 287 -31
rect 289 -41 295 -31
rect 297 -41 298 -31
rect 337 -41 338 -31
rect 340 -41 346 -31
rect 348 -41 349 -31
rect 369 -41 370 -31
rect 372 -41 378 -31
rect 380 -41 381 -31
rect 404 -41 405 -31
rect 407 -41 413 -31
rect 415 -41 416 -31
rect 444 -41 445 -31
rect 447 -41 453 -31
rect 455 -41 456 -31
rect 485 -41 486 -31
rect 488 -41 494 -31
rect 496 -41 497 -31
rect 519 -41 520 -31
rect 522 -41 528 -31
rect 530 -41 531 -31
rect 557 -41 558 -31
rect 560 -41 566 -31
rect 568 -41 569 -31
rect 595 -41 596 -31
rect 598 -41 604 -31
rect 606 -41 607 -31
rect 629 -41 630 -31
rect 632 -41 638 -31
rect 640 -41 641 -31
<< pdiffusion >>
rect -6 21 -5 41
rect -3 21 -2 41
rect 2 21 3 41
rect 5 21 6 41
rect 26 21 27 41
rect 29 21 30 41
rect 34 21 35 41
rect 37 21 38 41
rect 61 21 62 41
rect 64 21 65 41
rect 69 21 70 41
rect 72 21 73 41
rect 101 21 102 41
rect 104 21 105 41
rect 109 21 110 41
rect 112 21 113 41
rect 142 21 143 41
rect 145 21 146 41
rect 150 21 151 41
rect 153 21 154 41
rect 176 21 177 41
rect 179 21 180 41
rect 184 21 185 41
rect 187 21 188 41
rect 214 21 215 41
rect 217 21 218 41
rect 222 21 223 41
rect 225 21 226 41
rect 252 21 253 41
rect 255 21 256 41
rect 260 21 261 41
rect 263 21 264 41
rect 286 21 287 41
rect 289 21 290 41
rect 294 21 295 41
rect 297 21 298 41
rect 337 21 338 41
rect 340 21 341 41
rect 345 21 346 41
rect 348 21 349 41
rect 369 21 370 41
rect 372 21 373 41
rect 377 21 378 41
rect 380 21 381 41
rect 404 21 405 41
rect 407 21 408 41
rect 412 21 413 41
rect 415 21 416 41
rect 444 21 445 41
rect 447 21 448 41
rect 452 21 453 41
rect 455 21 456 41
rect 485 21 486 41
rect 488 21 489 41
rect 493 21 494 41
rect 496 21 497 41
rect 519 21 520 41
rect 522 21 523 41
rect 527 21 528 41
rect 530 21 531 41
rect 557 21 558 41
rect 560 21 561 41
rect 565 21 566 41
rect 568 21 569 41
rect 595 21 596 41
rect 598 21 599 41
rect 603 21 604 41
rect 606 21 607 41
rect 629 21 630 41
rect 632 21 633 41
rect 637 21 638 41
rect 640 21 641 41
<< ndcontact >>
rect -10 -41 -6 -31
rect 6 -41 10 -31
rect 22 -41 26 -31
rect 38 -41 42 -31
rect 57 -41 61 -31
rect 73 -41 77 -31
rect 97 -41 101 -31
rect 113 -41 117 -31
rect 138 -41 142 -31
rect 154 -41 158 -31
rect 172 -41 176 -31
rect 188 -41 192 -31
rect 210 -41 214 -31
rect 226 -41 230 -31
rect 248 -41 252 -31
rect 264 -41 268 -31
rect 282 -41 286 -31
rect 298 -41 302 -31
rect 333 -41 337 -31
rect 349 -41 353 -31
rect 365 -41 369 -31
rect 381 -41 385 -31
rect 400 -41 404 -31
rect 416 -41 420 -31
rect 440 -41 444 -31
rect 456 -41 460 -31
rect 481 -41 485 -31
rect 497 -41 501 -31
rect 515 -41 519 -31
rect 531 -41 535 -31
rect 553 -41 557 -31
rect 569 -41 573 -31
rect 591 -41 595 -31
rect 607 -41 611 -31
rect 625 -41 629 -31
rect 641 -41 645 -31
<< pdcontact >>
rect -10 21 -6 41
rect -2 21 2 41
rect 6 21 10 41
rect 22 21 26 41
rect 30 21 34 41
rect 38 21 42 41
rect 57 21 61 41
rect 65 21 69 41
rect 73 21 77 41
rect 97 21 101 41
rect 105 21 109 41
rect 113 21 117 41
rect 138 21 142 41
rect 146 21 150 41
rect 154 21 158 41
rect 172 21 176 41
rect 180 21 184 41
rect 188 21 192 41
rect 210 21 214 41
rect 218 21 222 41
rect 226 21 230 41
rect 248 21 252 41
rect 256 21 260 41
rect 264 21 268 41
rect 282 21 286 41
rect 290 21 294 41
rect 298 21 302 41
rect 333 21 337 41
rect 341 21 345 41
rect 349 21 353 41
rect 365 21 369 41
rect 373 21 377 41
rect 381 21 385 41
rect 400 21 404 41
rect 408 21 412 41
rect 416 21 420 41
rect 440 21 444 41
rect 448 21 452 41
rect 456 21 460 41
rect 481 21 485 41
rect 489 21 493 41
rect 497 21 501 41
rect 515 21 519 41
rect 523 21 527 41
rect 531 21 535 41
rect 553 21 557 41
rect 561 21 565 41
rect 569 21 573 41
rect 591 21 595 41
rect 599 21 603 41
rect 607 21 611 41
rect 625 21 629 41
rect 633 21 637 41
rect 641 21 645 41
<< psubstratepcontact >>
rect -9 -50 -5 -46
rect 5 -50 9 -46
rect 23 -50 27 -46
rect 37 -50 41 -46
rect 58 -50 62 -46
rect 72 -50 76 -46
rect 98 -50 102 -46
rect 112 -50 116 -46
rect 139 -50 143 -46
rect 153 -50 157 -46
rect 173 -50 177 -46
rect 187 -50 191 -46
rect 211 -50 215 -46
rect 225 -50 229 -46
rect 249 -50 253 -46
rect 263 -50 267 -46
rect 283 -50 287 -46
rect 297 -50 301 -46
rect 334 -50 338 -46
rect 348 -50 352 -46
rect 366 -50 370 -46
rect 380 -50 384 -46
rect 401 -50 405 -46
rect 415 -50 419 -46
rect 441 -50 445 -46
rect 455 -50 459 -46
rect 482 -50 486 -46
rect 496 -50 500 -46
rect 516 -50 520 -46
rect 530 -50 534 -46
rect 554 -50 558 -46
rect 568 -50 572 -46
rect 592 -50 596 -46
rect 606 -50 610 -46
rect 626 -50 630 -46
rect 640 -50 644 -46
<< nsubstratencontact >>
rect -9 46 -5 50
rect 5 46 9 50
rect 23 46 27 50
rect 37 46 41 50
rect 58 46 62 50
rect 72 46 76 50
rect 98 46 102 50
rect 112 46 116 50
rect 139 46 143 50
rect 153 46 157 50
rect 173 46 177 50
rect 187 46 191 50
rect 211 46 215 50
rect 225 46 229 50
rect 249 46 253 50
rect 263 46 267 50
rect 283 46 287 50
rect 297 46 301 50
rect 334 46 338 50
rect 348 46 352 50
rect 366 46 370 50
rect 380 46 384 50
rect 401 46 405 50
rect 415 46 419 50
rect 441 46 445 50
rect 455 46 459 50
rect 482 46 486 50
rect 496 46 500 50
rect 516 46 520 50
rect 530 46 534 50
rect 554 46 558 50
rect 568 46 572 50
rect 592 46 596 50
rect 606 46 610 50
rect 626 46 630 50
rect 640 46 644 50
<< polysilicon >>
rect -5 41 -3 44
rect 3 41 5 44
rect 27 41 29 44
rect 35 41 37 44
rect 62 41 64 44
rect 70 41 72 44
rect 102 41 104 44
rect 110 41 112 44
rect 143 41 145 44
rect 151 41 153 44
rect 177 41 179 44
rect 185 41 187 44
rect 215 41 217 44
rect 223 41 225 44
rect 253 41 255 44
rect 261 41 263 44
rect 287 41 289 44
rect 295 41 297 44
rect 338 41 340 44
rect 346 41 348 44
rect 370 41 372 44
rect 378 41 380 44
rect 405 41 407 44
rect 413 41 415 44
rect 445 41 447 44
rect 453 41 455 44
rect 486 41 488 44
rect 494 41 496 44
rect 520 41 522 44
rect 528 41 530 44
rect 558 41 560 44
rect 566 41 568 44
rect 596 41 598 44
rect 604 41 606 44
rect 630 41 632 44
rect 638 41 640 44
rect -5 16 -3 21
rect -7 12 -3 16
rect -5 -31 -3 12
rect 3 17 5 21
rect 3 13 7 17
rect 3 -31 5 13
rect 27 8 29 21
rect 24 4 29 8
rect 27 -31 29 4
rect 35 8 37 21
rect 62 17 64 21
rect 60 13 64 17
rect 35 4 39 8
rect 35 -31 37 4
rect 62 -31 64 13
rect 70 8 72 21
rect 102 17 104 21
rect 100 13 104 17
rect 70 4 74 8
rect 70 -31 72 4
rect 102 -31 104 13
rect 110 17 112 21
rect 143 17 145 21
rect 110 13 114 17
rect 141 13 145 17
rect 110 -31 112 13
rect 143 -31 145 13
rect 151 8 153 21
rect 177 17 179 21
rect 175 13 179 17
rect 151 4 155 8
rect 151 -31 153 4
rect 177 -31 179 13
rect 185 17 187 21
rect 215 17 217 21
rect 185 13 189 17
rect 213 13 217 17
rect 185 -31 187 13
rect 215 -31 217 13
rect 223 17 225 21
rect 253 17 255 21
rect 223 13 227 17
rect 251 13 255 17
rect 223 -31 225 13
rect 253 -31 255 13
rect 261 17 263 21
rect 287 17 289 21
rect 261 13 265 17
rect 285 13 289 17
rect 261 -31 263 13
rect 287 -31 289 13
rect 295 17 297 21
rect 295 13 299 17
rect 338 16 340 21
rect 295 -31 297 13
rect 336 12 340 16
rect 338 -31 340 12
rect 346 17 348 21
rect 346 13 350 17
rect 346 -31 348 13
rect 370 8 372 21
rect 367 4 372 8
rect 370 -31 372 4
rect 378 8 380 21
rect 405 17 407 21
rect 403 13 407 17
rect 378 4 382 8
rect 378 -31 380 4
rect 405 -31 407 13
rect 413 8 415 21
rect 445 17 447 21
rect 443 13 447 17
rect 413 4 417 8
rect 413 -31 415 4
rect 445 -31 447 13
rect 453 17 455 21
rect 486 17 488 21
rect 453 13 457 17
rect 484 13 488 17
rect 453 -31 455 13
rect 486 -31 488 13
rect 494 8 496 21
rect 520 17 522 21
rect 518 13 522 17
rect 494 4 498 8
rect 494 -31 496 4
rect 520 -31 522 13
rect 528 17 530 21
rect 558 17 560 21
rect 528 13 532 17
rect 556 13 560 17
rect 528 -31 530 13
rect 558 -31 560 13
rect 566 17 568 21
rect 596 17 598 21
rect 566 13 570 17
rect 594 13 598 17
rect 566 -31 568 13
rect 596 -31 598 13
rect 604 17 606 21
rect 630 17 632 21
rect 604 13 608 17
rect 628 13 632 17
rect 604 -31 606 13
rect 630 -31 632 13
rect 638 17 640 21
rect 638 13 642 17
rect 638 -31 640 13
rect -5 -44 -3 -41
rect 3 -44 5 -41
rect 27 -44 29 -41
rect 35 -44 37 -41
rect 62 -44 64 -41
rect 70 -44 72 -41
rect 102 -44 104 -41
rect 110 -44 112 -41
rect 143 -44 145 -41
rect 151 -44 153 -41
rect 177 -44 179 -41
rect 185 -44 187 -41
rect 215 -44 217 -41
rect 223 -44 225 -41
rect 253 -44 255 -41
rect 261 -44 263 -41
rect 287 -44 289 -41
rect 295 -44 297 -41
rect 338 -44 340 -41
rect 346 -44 348 -41
rect 370 -44 372 -41
rect 378 -44 380 -41
rect 405 -44 407 -41
rect 413 -44 415 -41
rect 445 -44 447 -41
rect 453 -44 455 -41
rect 486 -44 488 -41
rect 494 -44 496 -41
rect 520 -44 522 -41
rect 528 -44 530 -41
rect 558 -44 560 -41
rect 566 -44 568 -41
rect 596 -44 598 -41
rect 604 -44 606 -41
rect 630 -44 632 -41
rect 638 -44 640 -41
<< polycontact >>
rect -11 12 -7 16
rect 7 13 11 17
rect 20 4 24 8
rect 56 13 60 17
rect 39 4 43 8
rect 96 13 100 17
rect 74 4 78 8
rect 114 13 118 17
rect 137 13 141 17
rect 171 13 175 17
rect 155 4 159 8
rect 189 13 193 17
rect 209 13 213 17
rect 227 13 231 17
rect 247 13 251 17
rect 265 13 269 17
rect 281 13 285 17
rect 299 13 303 17
rect 332 12 336 16
rect 350 13 354 17
rect 363 4 367 8
rect 399 13 403 17
rect 382 4 386 8
rect 439 13 443 17
rect 417 4 421 8
rect 457 13 461 17
rect 480 13 484 17
rect 514 13 518 17
rect 498 4 502 8
rect 532 13 536 17
rect 552 13 556 17
rect 570 13 574 17
rect 590 13 594 17
rect 608 13 612 17
rect 624 13 628 17
rect 642 13 646 17
<< metal1 >>
rect -23 50 655 51
rect -23 46 -9 50
rect -5 46 5 50
rect 9 46 23 50
rect 27 46 37 50
rect 41 46 58 50
rect 62 46 72 50
rect 76 46 98 50
rect 102 46 112 50
rect 116 46 139 50
rect 143 46 153 50
rect 157 46 173 50
rect 177 46 187 50
rect 191 46 211 50
rect 215 46 225 50
rect 229 46 249 50
rect 253 46 263 50
rect 267 46 283 50
rect 287 46 297 50
rect 301 46 334 50
rect 338 46 348 50
rect 352 46 366 50
rect 370 46 380 50
rect 384 46 401 50
rect 405 46 415 50
rect 419 46 441 50
rect 445 46 455 50
rect 459 46 482 50
rect 486 46 496 50
rect 500 46 516 50
rect 520 46 530 50
rect 534 46 554 50
rect 558 46 568 50
rect 572 46 592 50
rect 596 46 606 50
rect 610 46 626 50
rect 630 46 640 50
rect 644 46 655 50
rect -23 45 655 46
rect -10 41 -6 45
rect 6 41 10 45
rect 22 41 26 45
rect 38 41 42 45
rect 57 41 61 45
rect 73 41 77 45
rect 97 41 101 45
rect 113 41 117 45
rect 138 41 142 45
rect 154 41 158 45
rect 172 41 176 45
rect 188 41 192 45
rect 210 41 214 45
rect 226 41 230 45
rect 248 41 252 45
rect 264 41 268 45
rect 282 41 286 45
rect 298 41 302 45
rect 333 41 337 45
rect 349 41 353 45
rect 365 41 369 45
rect 381 41 385 45
rect 400 41 404 45
rect 416 41 420 45
rect 440 41 444 45
rect 456 41 460 45
rect 481 41 485 45
rect 497 41 501 45
rect 515 41 519 45
rect 531 41 535 45
rect 553 41 557 45
rect 569 41 573 45
rect 591 41 595 45
rect 607 41 611 45
rect 625 41 629 45
rect 641 41 645 45
rect -17 16 -5 17
rect -17 12 -11 16
rect -7 12 -5 16
rect -17 11 -5 12
rect -2 0 2 21
rect 5 17 16 18
rect 5 13 7 17
rect 11 13 16 17
rect 14 4 20 8
rect 30 0 34 21
rect 50 17 60 18
rect 50 13 56 17
rect 50 12 60 13
rect 65 17 69 21
rect 95 17 100 18
rect 65 13 96 17
rect 100 13 102 17
rect 39 8 50 9
rect 43 4 50 8
rect 39 3 50 4
rect -2 -4 14 0
rect 6 -31 10 -4
rect 30 -4 42 0
rect 38 -15 42 -4
rect 45 -4 50 3
rect 65 0 69 13
rect 95 12 100 13
rect 74 8 85 9
rect 78 4 85 8
rect 74 3 85 4
rect 65 -4 77 0
rect 38 -20 54 -15
rect 38 -31 42 -20
rect 73 -31 77 -4
rect 80 -23 85 3
rect 105 0 109 21
rect 146 18 150 21
rect 114 17 125 18
rect 112 13 114 17
rect 118 13 125 17
rect 114 12 125 13
rect 120 5 125 12
rect 129 17 141 18
rect 146 17 175 18
rect 129 13 137 17
rect 141 13 143 17
rect 146 13 171 17
rect 175 13 177 17
rect 129 12 141 13
rect 146 12 175 13
rect 105 -4 117 0
rect 113 -24 117 -4
rect 129 -24 135 12
rect 146 0 150 12
rect 155 8 162 9
rect 159 4 162 8
rect 155 3 162 4
rect 180 0 184 21
rect 203 18 207 21
rect 189 17 199 18
rect 193 13 199 17
rect 203 17 213 18
rect 203 14 209 17
rect 189 12 199 13
rect 146 -4 158 0
rect 180 -4 192 0
rect 113 -29 130 -24
rect 154 -18 158 -4
rect 188 -14 192 -4
rect 195 -1 199 12
rect 207 13 209 14
rect 213 13 215 17
rect 154 -22 171 -18
rect 113 -31 117 -29
rect 154 -31 158 -22
rect 188 -19 195 -14
rect 188 -31 192 -19
rect 207 -23 213 13
rect 218 0 222 21
rect 240 18 244 21
rect 227 17 237 18
rect 231 13 237 17
rect 240 17 251 18
rect 240 14 247 17
rect 227 12 237 13
rect 245 13 247 14
rect 251 13 253 17
rect 245 12 251 13
rect 232 9 237 12
rect 256 9 260 21
rect 265 17 276 18
rect 269 13 276 17
rect 265 12 276 13
rect 256 5 263 9
rect 256 0 260 5
rect 218 -4 237 0
rect 212 -28 213 -23
rect 226 -5 237 -4
rect 256 -4 268 0
rect 226 -31 230 -5
rect 264 -31 268 -4
rect 271 -34 276 12
rect 280 17 285 18
rect 280 13 281 17
rect 285 13 287 17
rect 280 1 285 13
rect 290 0 294 21
rect 299 17 311 18
rect 297 13 299 17
rect 303 13 311 17
rect 299 12 311 13
rect 290 -4 302 0
rect 298 -31 302 -4
rect 306 -21 311 12
rect 326 16 338 17
rect 326 12 332 16
rect 336 12 338 16
rect 326 11 338 12
rect 341 0 345 21
rect 348 17 359 18
rect 348 13 350 17
rect 354 13 359 17
rect 357 8 367 9
rect 357 4 363 8
rect 373 0 377 21
rect 393 17 403 18
rect 393 13 399 17
rect 393 12 403 13
rect 408 17 412 21
rect 438 17 443 18
rect 408 13 439 17
rect 443 13 445 17
rect 382 8 393 9
rect 386 4 393 8
rect 382 3 393 4
rect 341 -4 357 0
rect 349 -31 353 -4
rect 373 -4 385 0
rect 381 -15 385 -4
rect 388 -4 393 3
rect 408 0 412 13
rect 438 12 443 13
rect 417 8 428 9
rect 421 4 428 8
rect 417 3 428 4
rect 408 -4 420 0
rect 381 -20 397 -15
rect 381 -31 385 -20
rect 416 -31 420 -4
rect 423 -23 428 3
rect 448 0 452 21
rect 489 18 493 21
rect 457 17 468 18
rect 455 13 457 17
rect 461 13 468 17
rect 457 12 468 13
rect 463 5 468 12
rect 472 17 484 18
rect 489 17 518 18
rect 472 13 480 17
rect 484 13 486 17
rect 489 13 514 17
rect 518 13 520 17
rect 472 12 484 13
rect 489 12 518 13
rect 448 -4 460 0
rect 456 -24 460 -4
rect 472 -24 478 12
rect 489 0 493 12
rect 498 8 505 9
rect 502 4 505 8
rect 498 3 505 4
rect 523 0 527 21
rect 546 18 550 21
rect 532 17 542 18
rect 536 13 542 17
rect 546 17 556 18
rect 546 14 552 17
rect 532 12 542 13
rect 489 -4 501 0
rect 523 -4 535 0
rect 456 -29 473 -24
rect 497 -18 501 -4
rect 531 -14 535 -4
rect 538 -1 542 12
rect 550 13 552 14
rect 556 13 558 17
rect 497 -22 514 -18
rect 456 -31 460 -29
rect 497 -31 501 -22
rect 531 -19 538 -14
rect 531 -31 535 -19
rect 550 -23 556 13
rect 561 0 565 21
rect 583 18 587 21
rect 570 17 580 18
rect 574 13 580 17
rect 583 17 594 18
rect 583 14 590 17
rect 570 12 580 13
rect 588 13 590 14
rect 594 13 596 17
rect 588 12 594 13
rect 575 9 580 12
rect 599 0 603 21
rect 608 17 619 18
rect 612 13 619 17
rect 608 12 619 13
rect 561 -4 580 0
rect 555 -28 556 -23
rect 569 -5 580 -4
rect 599 -4 611 0
rect 569 -31 573 -5
rect 607 -31 611 -4
rect 614 -34 619 12
rect 623 17 628 18
rect 623 13 624 17
rect 628 13 630 17
rect 623 1 628 13
rect 633 0 637 21
rect 642 17 654 18
rect 640 13 642 17
rect 646 13 654 17
rect 642 12 654 13
rect 633 -4 645 0
rect 641 -31 645 -4
rect 649 -21 654 12
rect -10 -45 -6 -41
rect 22 -45 26 -41
rect 57 -45 61 -41
rect 97 -45 101 -41
rect 138 -45 142 -41
rect 172 -45 176 -41
rect 210 -45 214 -41
rect 248 -45 252 -41
rect 282 -45 286 -41
rect 333 -45 337 -41
rect 365 -45 369 -41
rect 400 -45 404 -41
rect 440 -45 444 -41
rect 481 -45 485 -41
rect 515 -45 519 -41
rect 553 -45 557 -41
rect 591 -45 595 -41
rect 625 -45 629 -41
rect -23 -46 655 -45
rect -23 -50 -9 -46
rect -5 -50 5 -46
rect 9 -50 23 -46
rect 27 -50 37 -46
rect 41 -50 58 -46
rect 62 -50 72 -46
rect 76 -50 98 -46
rect 102 -50 112 -46
rect 116 -50 139 -46
rect 143 -50 153 -46
rect 157 -50 173 -46
rect 177 -50 187 -46
rect 191 -50 211 -46
rect 215 -50 225 -46
rect 229 -50 249 -46
rect 253 -50 263 -46
rect 267 -50 283 -46
rect 287 -50 297 -46
rect 301 -50 334 -46
rect 338 -50 348 -46
rect 352 -50 366 -46
rect 370 -50 380 -46
rect 384 -50 401 -46
rect 405 -50 415 -46
rect 419 -50 441 -46
rect 445 -50 455 -46
rect 459 -50 482 -46
rect 486 -50 496 -46
rect 500 -50 516 -46
rect 520 -50 530 -46
rect 534 -50 554 -46
rect 558 -50 568 -46
rect 572 -50 592 -46
rect 596 -50 606 -46
rect 610 -50 626 -46
rect 630 -50 640 -46
rect 644 -50 655 -46
rect -23 -51 655 -50
<< m2contact >>
rect 202 21 207 26
rect 239 21 244 26
rect 545 21 550 26
rect 582 21 587 26
rect -23 11 -17 17
rect 16 13 21 18
rect 8 4 14 9
rect 44 12 50 18
rect 14 -5 19 0
rect 45 -9 50 -4
rect 54 -19 59 -14
rect 120 0 125 5
rect 80 -28 85 -23
rect 162 3 167 9
rect 130 -29 135 -24
rect 195 -6 200 -1
rect 171 -23 176 -18
rect 195 -19 200 -14
rect 232 4 237 9
rect 263 4 268 9
rect 207 -28 212 -23
rect 237 -5 242 0
rect 280 -4 285 1
rect 320 11 326 17
rect 359 13 364 18
rect 351 4 357 9
rect 387 12 393 18
rect 306 -26 311 -21
rect 357 -5 362 0
rect 388 -9 393 -4
rect 397 -19 402 -14
rect 463 0 468 5
rect 423 -28 428 -23
rect 505 4 510 9
rect 473 -29 478 -24
rect 538 -6 543 -1
rect 514 -23 519 -18
rect 538 -19 543 -14
rect 575 4 580 9
rect 550 -28 555 -23
rect 580 -5 585 0
rect 271 -39 276 -34
rect 623 -4 628 1
rect 649 -26 654 -21
rect 614 -39 619 -34
<< metal2 >>
rect 312 37 509 41
rect 207 21 239 26
rect 21 13 44 18
rect -23 9 -17 11
rect 312 9 316 37
rect -23 3 8 9
rect 167 4 232 9
rect 268 5 316 9
rect 364 12 387 18
rect 320 9 326 11
rect 505 9 509 37
rect 550 21 582 26
rect 320 3 351 9
rect 14 -10 19 -5
rect 45 -10 50 -9
rect 14 -15 50 -10
rect 120 -14 125 0
rect 45 -23 50 -15
rect 59 -19 125 -14
rect 162 -6 195 -1
rect 242 -4 280 0
rect 510 4 575 9
rect 45 -28 80 -23
rect 85 -28 125 -23
rect 162 -24 167 -6
rect 357 -10 362 -5
rect 388 -10 393 -9
rect 120 -34 125 -28
rect 135 -29 167 -24
rect 200 -19 244 -14
rect 357 -15 393 -10
rect 463 -14 468 0
rect 239 -22 244 -19
rect 171 -28 207 -23
rect 239 -26 306 -22
rect 388 -23 393 -15
rect 402 -19 468 -14
rect 505 -6 538 -1
rect 585 -4 623 0
rect 388 -28 423 -23
rect 428 -28 468 -23
rect 505 -24 510 -6
rect 463 -34 468 -28
rect 478 -29 510 -24
rect 543 -19 587 -14
rect 582 -22 587 -19
rect 514 -28 550 -23
rect 582 -26 649 -22
rect 120 -39 271 -34
rect 463 -39 614 -34
<< labels >>
rlabel metal1 -1 -49 -1 -49 1 GND
rlabel metal1 609 -7 609 -7 1 COUT
rlabel metal1 0 48 0 48 5 VDD
rlabel polysilicon 152 6 152 6 1 C
rlabel polysilicon -4 11 -4 11 1 A
rlabel polysilicon 4 11 4 11 1 B
rlabel metal1 300 -7 300 -7 1 Y
rlabel polysilicon 339 11 339 11 1 D
rlabel polysilicon 347 11 347 11 1 E
rlabel metal1 643 -7 643 -7 1 Z
<< end >>
